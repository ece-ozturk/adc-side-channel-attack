** Simulation of synthesized D flip-flop circuit with NGSpice

** Include necessary library and synthesized model file
.lib "/foss/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.include "/foss/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice"
.include dff_corrected_synth.model

** Instantiate the D flip-flop module
Xdff clk rst d q vss vss vdd vdd dff

** Define power supply
.param vss=0
Vvss vss 0 {vss}

** Define power supply
.param vdd=1.8
Vvdd vdd 0 {vdd}

** Clock signal: 2 MHz, 50% duty cycle
Vclk clk 0 pulse 0 {vdd} 200n 10n 10n 1u 2u

** Reset signal: Pulse for the first few cycles to initialize
Vrst rst 0 pulse {vdd} 500n 0 5n 5n 10u 15u

** Enable signal: Enable after reset
** Ven en 0 pulse 0 {vdd} 1u 5n 5n 500n 3u

** Data input: Toggles every 2 µs
Vd d 0 pulse 0 {vdd} 1u 5n 5n 2.5u 6u

** Simulation control
.control
    tran 100n 40u 0 1n
    plot (clk) (rst) (d) (q)
.endc
.END
